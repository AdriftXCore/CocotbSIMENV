package dff_pkg;

parameter TEST_PKG = 32'h20251121;
parameter TEST_PKG1 = 32'h5a5aa5a5;

endpackage